`timescale 1ns/1ps
module tb_int_receiver ();
    
endmodule