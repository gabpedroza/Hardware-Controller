`timescale 1ns/1ps
module send_receive_test();

    

endmodule